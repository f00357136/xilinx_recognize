`include "define.v"
module WRA_Top
// ----------------------------------------------------------------------------
// Port declarations
// ----------------------------------------------------------------------------
(input  wire [`WRAInAddrWidth-1:0] a,
 input  wire clk,
 input  wire rst,
 input  wire stride_op,
 input  wire kernelsize_op,
 input  wire inputbstart_op,
 input  wire poolingen_op,
 input  wire padding_op,
 input  wire [8:0] numslideH_op, //max=510 大小�?1024，min=3 大小�?8,  多个输入通道组成 
 input  wire [4:0] numslideV_op, //max=31
 input  wire [4:0] numswitchH_op, //横向窗口滑动通道转换距离
 input  wire [4:0] NInch_D_PInch_op, //max=512/16=32
 input  wire [4:0] NOuch_D_POuch_op, //max=512/16=32
 input  wire [7:0] cellnum_op,
 input  wire [7:0] linenum_op,
 input  wire [1:0] fixpoint_op,
 input  wire relu_op,
 input  wire [`AyInFIFOWidth-1:0] d_ram,
 input  wire we,
 input  wire we_Gt,
 input  wire [`AyFiFIFOWidth-1:0] d_Gt,
 input  wire [`FiBufferSize-1:0]  a_GtOutside,
 output wire Layer_Finish,
 output wire [`WRAOutDataWidth-1:0]WRA_FeatureData
 );
 
/*-----------------------------------------------------------------------------------------------------------------------*/
/*-----------------------------------------------------------------------------------------------------------------------*/
wire [3:0] current_state;
wire [3:0] current_state_d;
wire [3:0] current_state_4d;
wire [3:0] current_state_5d;

wire [`FiBufferSize-1:0] a_Gt, a_Gt1, a_Gt2;
wire [`InBuOutDaWidth-1:0] inputb_spo;
wire [`NumBuLine-1:0]ex_we, ex_we_padding; 
wire [7:0] ex_addr;	
wire [`InBuInDaWidthMax-1:0] ex_d1, ex_d2;
assign a_Gt1=a_GtOutside;
assign a_Gt=(we_Gt==1)?a_Gt1:a_Gt2;

Input_Buffer Input_Buffer0(
    .a(a),                              //Inout Buffer READ address, for capturing data from Inout Buffer to AHB read_data
									    //Generated by AHB reg_haddr from WAR_SLAVE
    .d(d_ram),							//Inout Buffer input data, 128 bit width, can be set according by Feature FIFO output 
										//data width
    .we(we),                            //Inout Buffer input data write enable
    .clk(clk), 
    .inputb_spo(inputb_spo),            //Multiple-channels output data
    .rst(rst), 
    .stride_op(stride_op),      
    .kernelsize_op(kernelsize_op), 
    .numslideH_op(numslideH_op),
    .numslideV_op(numslideV_op),
    .BtInB_Save_Done(BtInB_Save_Done),  //Represent all the TILES DATA needed in one 4-ROWS computation of one layer has been
										//transformed (or not) and saved in BtInB_Buffer 
    .en_accord_inputbstart(en_accord_inputbstart), 
										//Enable BtInB transformation and BtInB_Buffer saving 
    .ex_we(ex_we),                      //Exchange enable when output data restores in Inout Buffer
    .ex_addr(ex_addr),                  //Exchange address when output data restores in Inout Buffer
    .ex_d1(ex_d1),                      //First  row Exchange data
    .ex_d2(ex_d2), 						//Second row Exchange data
    .current_state(current_state),      
    .Channel_Switch_Done_6d(Channel_Switch_Done_6d), 
										//A pulse indicates one 4-ROWS computation and restoring of one layer has been done 
    .Layer_Finish(Layer_Finish),        //A pulse indicates one layer of CNN model has been done
    .numswitchH_op(numswitchH_op), 
    .poolingen_op(poolingen_op), 
    .cellnum_op(cellnum_op),            //Represent how much feature data need to be initiated in one "Buffer_Grain_16_32_32bit"
										//model
    .linenum_op(linenum_op),            //Represent how many line data need to be initiated in Inout Buffer
    .ex_we_padding(ex_we_padding),      //Padding enable while BtInB Transformation is running
    .WRA_FeatureData(WRA_FeatureData)   //Inout Buffer READ data, provided to AHB read_data
);

wire [`InTrOutDaWidth-1 :0] output16_8bit1;
wire [`InTrOutDaWidth-1 :0] output16_8bit2;
wire [`InTrOutDaWidth-1 :0] output16_8bit3;
wire [`InTrOutDaWidth-1 :0] output16_8bit4;

Input_Trans Input_Trans1 (				//Cut according to input channel
    .input16_8bit(inputb_spo[127 :0	  ]),									
    .clk(clk), 
    .rst(rst), 
    .output16_8bit(output16_8bit1),     
    .fixpoint_op(fixpoint_op)
);

Input_Trans Input_Trans2 (
    .input16_8bit(inputb_spo[255 :128 ]), 
    .clk(clk), 
    .rst(rst), 
    .output16_8bit(output16_8bit2), 
    .fixpoint_op(fixpoint_op)
);

Input_Trans Input_Trans3 (
    .input16_8bit(inputb_spo[383 :256 ]), 
    .clk(clk), 
    .rst(rst), 
    .output16_8bit(output16_8bit3), 
    .fixpoint_op(fixpoint_op)
);

Input_Trans Input_Trans4 (
    .input16_8bit(inputb_spo[511 :384 ]), 
    .clk(clk), 
    .rst(rst), 
    .output16_8bit(output16_8bit4), 
    .fixpoint_op(fixpoint_op)
);

wire [`BtBuDaWidth-1:0] BtInB_spo;
assign BtInB_spo={output16_8bit4,
				  output16_8bit3,
				  output16_8bit2,
				  output16_8bit1};	
			  
wire [`BtBuDaWidth-1:0] BtInB_RAMspo;
wire [3:0] a_Bt;

BtInB_Buffer BtInB_Buffer0(
    .BtInB_spo(BtInB_spo),
    .inputb_spo(inputb_spo),
    .a_Bt(a_Bt),
    .clk(clk),
    .we_Bt(we_Bt),
    .spo(BtInB_RAMspo),
    .kernelsize_op(kernelsize_op)
);

wire [`GtBuDaWidth-1:0] GFGt_RAMspo;

GFGt_Ram GFGt_Ram0(
	.clk(clk), 
	.we(we_Gt), 
	.a(a_Gt), 
	.d(d_Gt), 
	.spo(GFGt_RAMspo)
);  

wire [`GtInDSPWidth-1:0]GFGt1,GFGt2,GFGt3,GFGt4;

assign GFGt1=GFGt_RAMspo[511 :0   ];//Cut according to output channel
assign GFGt2=GFGt_RAMspo[1023:512 ];
assign GFGt3=GFGt_RAMspo[1535:1024];
assign GFGt4=GFGt_RAMspo[2047:1536];

wire [`DSPOutWidthA-1:0]UpV1,UpV2,UpV3,UpV4;

DSP16_16 DSP16_1 ( //Cut according to input channel
	.clk(clk), 
	.inputa(BtInB_RAMspo), 
	.inputb(GFGt1), 
	.outputp(UpV1),
	.fixpoint_op(fixpoint_op)
);

DSP16_16 DSP16_2 ( //Cut according to input channel
	.clk(clk), 
	.inputa(BtInB_RAMspo), 
	.inputb(GFGt2), 
	.outputp(UpV2),
	.fixpoint_op(fixpoint_op)
);

DSP16_16 DSP16_3 ( //Cut according to input channel
	.clk(clk), 
	.inputa(BtInB_RAMspo), 
	.inputb(GFGt3), 
	.outputp(UpV3),
	.fixpoint_op(fixpoint_op)
);
//20190925 11:38�Ķ�
DSP16_16 DSP16_4 ( //Cut according to input channel
	.clk(clk), 
	.inputa(BtInB_RAMspo), 
	.inputb(GFGt4), 
	.outputp(UpV4),
	.fixpoint_op(fixpoint_op)
);

wire [`ChAcOutWidthA-1:0] UpV_Accumu1_16_1,UpV_Accumu1_16_2,UpV_Accumu1_16_3,UpV_Accumu1_16_4;

Channel_Accumu1_16 Channel_Accumu1_16_1 (//Cut according to input channel
	.clk(clk), 
	.rst(rst), 
	.UpV(UpV1), 
	.UpV_Accumu1_16(UpV_Accumu1_16_1)
);
 
Channel_Accumu1_16 Channel_Accumu1_16_2 (
	.clk(clk), 
	.rst(rst), 
	.UpV(UpV2), 
	.UpV_Accumu1_16(UpV_Accumu1_16_2)
);

Channel_Accumu1_16 Channel_Accumu1_16_3 (
	.clk(clk), 
	.rst(rst), 
	.UpV(UpV3), 
	.UpV_Accumu1_16(UpV_Accumu1_16_3)
);
//20190925 11:38�Ķ�
Channel_Accumu1_16 Channel_Accumu1_16_4 (
	.clk(clk), 
	.rst(rst), 
	.UpV(UpV4), 
	.UpV_Accumu1_16(UpV_Accumu1_16_4)
); 

wire [`ChAcNOutWidthA-1:0] UpV_Accumu1_N_1,UpV_Accumu1_N_2,UpV_Accumu1_N_3,UpV_Accumu1_N_4;

Channel_Accumulator Channel_Accumulator1 ( //Cut according to output channel
	.clk(clk), 
	.rst(rst), 
	.current_state_5d(current_state_5d), 
	.UpV_Accumu1_16(UpV_Accumu1_16_1), 
	.UpV_Accumu1_N(UpV_Accumu1_N_1),
	.NInch_D_PInch_op(NInch_D_PInch_op),
	.UpV_Accumu1_N_en(UpV_Accumu1_N_en),
	.current_state_4d(current_state_4d)
);

Channel_Accumulator Channel_Accumulator2 (
	.clk(clk), 
	.rst(rst), 
	.current_state_5d(current_state_5d), 
	.UpV_Accumu1_16(UpV_Accumu1_16_2), 
	.UpV_Accumu1_N(UpV_Accumu1_N_2),
	.NInch_D_PInch_op(NInch_D_PInch_op),
	.current_state_4d(current_state_4d)
);

Channel_Accumulator Channel_Accumulator3 (
	.clk(clk), 
	.rst(rst), 
	.current_state_5d(current_state_5d), 
	.UpV_Accumu1_16(UpV_Accumu1_16_3), 
	.UpV_Accumu1_N(UpV_Accumu1_N_3),
	.NInch_D_PInch_op(NInch_D_PInch_op),
	.current_state_4d(current_state_4d)
);
//20190925 11:38�Ķ�
Channel_Accumulator Channel_Accumulator4 (
	.clk(clk), 
	.rst(rst), 
	.current_state_5d(current_state_5d), 
	.UpV_Accumu1_16(UpV_Accumu1_16_4), 
	.UpV_Accumu1_N(UpV_Accumu1_N_4),
	.NInch_D_PInch_op(NInch_D_PInch_op),
	.current_state_4d(current_state_4d)
);

wire [`OuTrDaWidth-1:0] AtUVA_B1_1; wire [`OuTrDaWidth-1:0] AtUVA_B2_1;
wire [`OuTrDaWidth-1:0] AtUVA_B1_2; wire [`OuTrDaWidth-1:0] AtUVA_B2_2;
wire [`OuTrDaWidth-1:0] AtUVA_B1_3; wire [`OuTrDaWidth-1:0] AtUVA_B2_3;
wire [`OuTrDaWidth-1:0] AtUVA_B1_4; wire [`OuTrDaWidth-1:0] AtUVA_B2_4;  //OuTrDaWidth=32
 
Output_Trans Output_Trans1 ( //Cut according to output channel
	.clk(clk) , 
	.UpV(UpV_Accumu1_N_1) , 
	.AtUVA_B1(AtUVA_B1_1) , 
	.AtUVA_B2(AtUVA_B2_1) , 
	.poolingen_op(poolingen_op) , 
	.kernelsize_op(kernelsize_op), 
	.relu_op(relu_op)
);

Output_Trans Output_Trans2 (
	.clk(clk) , 
	.UpV(UpV_Accumu1_N_2) , 
	.AtUVA_B1(AtUVA_B1_2) , 
	.AtUVA_B2(AtUVA_B2_2) , 
	.poolingen_op(poolingen_op) , 
	.kernelsize_op(kernelsize_op), 
	.relu_op(relu_op)
);

Output_Trans Output_Trans3 (
	.clk(clk) , 
	.UpV(UpV_Accumu1_N_3) , 
	.AtUVA_B1(AtUVA_B1_3) , 
	.AtUVA_B2(AtUVA_B2_3) , 
	.poolingen_op(poolingen_op) , 
	.kernelsize_op(kernelsize_op), 
	.relu_op(relu_op)
);
//20190925 11:38�Ķ�
Output_Trans Output_Trans4 (
	.clk(clk) , 
	.UpV(UpV_Accumu1_N_4) , 
	.AtUVA_B1(AtUVA_B1_4) , 
	.AtUVA_B2(AtUVA_B2_4) , 
	.poolingen_op(poolingen_op) , 
	.kernelsize_op(kernelsize_op), 
	.relu_op(relu_op)
);
//20190925 11:38�Ķ�
assign ex_d1=
{AtUVA_B1_4, AtUVA_B1_3, AtUVA_B1_2, AtUVA_B1_1};
assign ex_d2=
{AtUVA_B2_4, AtUVA_B2_3, AtUVA_B2_2, AtUVA_B2_1};

//assign ex_d1=
//{32'b0, AtUVA_B1_3, AtUVA_B1_2, AtUVA_B1_1};
//assign ex_d2=
//{32'b0, AtUVA_B2_3, AtUVA_B2_2, AtUVA_B2_1};


Buffer_Exchanger Buffer_Exchanger0(
	.clk(clk), 
	.rst(rst), 
	.current_state_5d(current_state_5d), 
	.UpV_Accumu1_N_en(UpV_Accumu1_N_en), 
	.ex_we(ex_we), 
	.ex_addr(ex_addr), 
	.numslideH_op(numslideH_op),
	.numswitchH_op(numswitchH_op), 
	.NInch_D_PInch_op(NInch_D_PInch_op), 
	.NOuch_D_POuch_op(NOuch_D_POuch_op), 
	.Layer_Finish(Layer_Finish), 
	.Channel_Switch_Done_6d(Channel_Switch_Done_6d), 
	.poolingen_op(poolingen_op),
	.inputbstart_op(inputbstart_op), 
	.en_accord_inputbstart(en_accord_inputbstart), 
	.ex_we_padding(ex_we_padding), 
	.padding_op(padding_op), 
	.kernelsize_op(kernelsize_op)
);

WRA_ctl WRA_ctl0(
	.clk(clk), 
	.rst(rst), 
	.BtInB_Save_Done(BtInB_Save_Done), 
	.Layer_Finish(Layer_Finish), 
	.Channel_Switch_Done_6d(Channel_Switch_Done_6d), 
	.inputbstart_op(inputbstart_op), 
	.numslideH_op(numslideH_op), 
	.numswitchH_op(numswitchH_op), 
	.numslideV_op(numslideV_op), 
	.NInch_D_PInch_op(NInch_D_PInch_op), 
	.NOuch_D_POuch_op(NOuch_D_POuch_op), 
	.en_accord_inputbstart(en_accord_inputbstart), 
	.we_Bt(we_Bt), 
	.a_Bt(a_Bt), 
	.a_Gt(a_Gt2), 
	.current_state_5d(current_state_5d), 
	.current_state(current_state), 
	.current_state_d(current_state_d), 
	.current_state_4d(current_state_4d)
);		

endmodule














